module CLK_GATING (
input 										CLK,
input 										EN,
output 										GATED_CLK
);

////////////////////////////////////////////////////////
///////////////// INTERNAL SIGNALS ///////////////////// 
////////////////////////////////////////////////////////

reg								 			o_latch;

////////////////////////////////////////////////////////
///////////////////// CLOCK GATING ///////////////////// 
////////////////////////////////////////////////////////

always @ (CLK or EN) begin
	if (!CLK)
	o_latch = EN;
end 

assign GATED_CLK = o_latch & CLK;

endmodule
